library IEEE;
use IEEE.std_logic_1164.all;

entity registerMEM_WB is

 generic(N : integer := 32); 

  port(i_CLK          : in std_logic;     -- Clock input
       i_RST          : in std_logic;     -- Reset input
       i_WE           : in std_logic;     -- Write enable input

       i_MemtoReg     : in std_logic; 
       i_regWrite     : in std_logic; 
       i_JumpLink     : in std_logic; 
       i_halt         : in std_logic; 
       i_regDst       : in std_logic;
       i_PCplus4      : in std_logic_vector(N-1 downto 0);
       i_DMEM         : in std_logic_vector(N-1 downto 0);
       i_ALU          : in std_logic_vector(N-1 downto 0);
       i_reg_addr     : in std_logic_vector(4 downto 0);

       o_MemtoReg     : out std_logic; 
       o_regWrite     : out std_logic; 
       o_JumpLink     : out std_logic; 
       o_halt         : out std_logic; 
       o_regDst       : out std_logic;
       o_PCplus4      : out std_logic_vector(N-1 downto 0);
       o_DMEM         : out std_logic_vector(N-1 downto 0);
       o_ALU          : out std_logic_vector(N-1 downto 0);
       o_reg_addr     : out std_logic_vector(4 downto 0));


end registerMEM_WB;


architecture behavioral of registerMEM_WB is

component n_bit_reg is
   generic(N : integer := 32);
  port(i_CLK        : in std_logic;   
       i_RST        : in std_logic;   
       i_WE         : in std_logic;  
       i_D          : in std_logic_vector(N-1 downto 0);
       o_Q          : out std_logic_vector(N-1 downto 0));
  end component;


component dffg is
  port(i_CLK        : in std_logic;     -- Clock input
       i_RST        : in std_logic;     -- Reset input
       i_WE         : in std_logic;     -- Write enable input
       i_D          : in std_logic;     -- Data value input
       o_Q          : out std_logic);   -- Data value output
  end component;


begin

    Csignal_reg_Dst: dffg         
      port map(i_D            => i_regDst,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_regDst); 

    Csignal_MemtoReg: dffg 
      port map(i_D            => i_MemtoReg,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_MemtoReg);    
  

    Csignal_regWrite: dffg 
      port map(i_D            => i_regWrite,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_regWrite);      

    Csignal_JumpLink: dffg 
      port map(i_D            => i_JumpLink,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_JumpLink);     

    Csignal_halt: dffg 
      port map(i_D            => i_halt,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_halt);    

    PCplus4: n_bit_reg 
      port map(i_D            => i_PCplus4,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_PCplus4);     

    DMEM: n_bit_reg 
      port map(i_D            => i_DMEM,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_DMEM);  

    ALU: n_bit_reg 
      port map(i_D            => i_ALU,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_ALU);   

    reg_addr: n_bit_reg 
  generic map(N => 5) 
      port map(i_D            => i_reg_addr,
               i_CLK          => i_CLK,
               i_RST          => i_RST,
               i_WE           => i_WE,
               o_Q            => o_reg_addr);      
 


  
end behavioral;
