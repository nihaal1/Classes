// Copyright (C) 2020  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 20.1.1 Build 720 11/11/2020 SJ Standard Edition"
// CREATED		"Wed Apr 27 17:39:25 2022"

module \2_to_4_decoder (
	w0,
	w1,
	En,
	y0,
	y1,
	y2,
	y3
);


input wire	w0;
input wire	w1;
input wire	En;
output wire	y0;
output wire	y1;
output wire	y2;
output wire	y3;

wire	SYNTHESIZED_WIRE_4;
wire	SYNTHESIZED_WIRE_5;




assign	y0 = SYNTHESIZED_WIRE_4 & En & SYNTHESIZED_WIRE_5;

assign	y1 = w0 & En & SYNTHESIZED_WIRE_5;

assign	y2 = w1 & En & SYNTHESIZED_WIRE_4;

assign	SYNTHESIZED_WIRE_4 =  ~w0;

assign	SYNTHESIZED_WIRE_5 =  ~w1;

assign	y3 = w0 & En & w1;


endmodule
